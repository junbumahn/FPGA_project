module de_serializer (
    input        i_pixclk       ,
    input        i_tmdsclk      ,
    input        i_serial_data  ,
    output [9:0] o_encoded_data ,
    
    
);
    
endmodule